library verilog;
use verilog.vl_types.all;
entity lab3_mm_interconnect_0 is
    port(
        hps_0_h2f_lw_axi_master_awid: in     vl_logic_vector(11 downto 0);
        hps_0_h2f_lw_axi_master_awaddr: in     vl_logic_vector(20 downto 0);
        hps_0_h2f_lw_axi_master_awlen: in     vl_logic_vector(3 downto 0);
        hps_0_h2f_lw_axi_master_awsize: in     vl_logic_vector(2 downto 0);
        hps_0_h2f_lw_axi_master_awburst: in     vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_awlock: in     vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_awcache: in     vl_logic_vector(3 downto 0);
        hps_0_h2f_lw_axi_master_awprot: in     vl_logic_vector(2 downto 0);
        hps_0_h2f_lw_axi_master_awvalid: in     vl_logic;
        hps_0_h2f_lw_axi_master_awready: out    vl_logic;
        hps_0_h2f_lw_axi_master_wid: in     vl_logic_vector(11 downto 0);
        hps_0_h2f_lw_axi_master_wdata: in     vl_logic_vector(31 downto 0);
        hps_0_h2f_lw_axi_master_wstrb: in     vl_logic_vector(3 downto 0);
        hps_0_h2f_lw_axi_master_wlast: in     vl_logic;
        hps_0_h2f_lw_axi_master_wvalid: in     vl_logic;
        hps_0_h2f_lw_axi_master_wready: out    vl_logic;
        hps_0_h2f_lw_axi_master_bid: out    vl_logic_vector(11 downto 0);
        hps_0_h2f_lw_axi_master_bresp: out    vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_bvalid: out    vl_logic;
        hps_0_h2f_lw_axi_master_bready: in     vl_logic;
        hps_0_h2f_lw_axi_master_arid: in     vl_logic_vector(11 downto 0);
        hps_0_h2f_lw_axi_master_araddr: in     vl_logic_vector(20 downto 0);
        hps_0_h2f_lw_axi_master_arlen: in     vl_logic_vector(3 downto 0);
        hps_0_h2f_lw_axi_master_arsize: in     vl_logic_vector(2 downto 0);
        hps_0_h2f_lw_axi_master_arburst: in     vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_arlock: in     vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_arcache: in     vl_logic_vector(3 downto 0);
        hps_0_h2f_lw_axi_master_arprot: in     vl_logic_vector(2 downto 0);
        hps_0_h2f_lw_axi_master_arvalid: in     vl_logic;
        hps_0_h2f_lw_axi_master_arready: out    vl_logic;
        hps_0_h2f_lw_axi_master_rid: out    vl_logic_vector(11 downto 0);
        hps_0_h2f_lw_axi_master_rdata: out    vl_logic_vector(31 downto 0);
        hps_0_h2f_lw_axi_master_rresp: out    vl_logic_vector(1 downto 0);
        hps_0_h2f_lw_axi_master_rlast: out    vl_logic;
        hps_0_h2f_lw_axi_master_rvalid: out    vl_logic;
        hps_0_h2f_lw_axi_master_rready: in     vl_logic;
        clk_0_clk_clk   : in     vl_logic;
        hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset: in     vl_logic;
        master_0_clk_reset_reset_bridge_in_reset_reset: in     vl_logic;
        vga_led_0_reset_sink_reset_bridge_in_reset_reset: in     vl_logic;
        master_0_master_address: in     vl_logic_vector(31 downto 0);
        master_0_master_waitrequest: out    vl_logic;
        master_0_master_byteenable: in     vl_logic_vector(3 downto 0);
        master_0_master_read: in     vl_logic;
        master_0_master_readdata: out    vl_logic_vector(31 downto 0);
        master_0_master_readdatavalid: out    vl_logic;
        master_0_master_write: in     vl_logic;
        master_0_master_writedata: in     vl_logic_vector(31 downto 0);
        vga_led_0_avalon_slave_0_address: out    vl_logic_vector(2 downto 0);
        vga_led_0_avalon_slave_0_write: out    vl_logic;
        vga_led_0_avalon_slave_0_writedata: out    vl_logic_vector(7 downto 0);
        vga_led_0_avalon_slave_0_chipselect: out    vl_logic
    );
end lab3_mm_interconnect_0;
