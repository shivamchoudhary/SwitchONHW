module RamScheduler(input clk,
        input in_ram1,in_ram2,in_ram3
);
        
        function logic set_rd(logic [31:0] data, logic[1:0] in, logic [1:0]size)


        always_ff @(posedge clk)
                in_rd_ram1 = 

