library verilog;
use verilog.vl_types.all;
entity lab3_hps_0_hps_io is
    port(
        mem_a           : out    vl_logic_vector(14 downto 0);
        mem_ba          : out    vl_logic_vector(2 downto 0);
        mem_ck          : out    vl_logic;
        mem_ck_n        : out    vl_logic;
        mem_cke         : out    vl_logic;
        mem_cs_n        : out    vl_logic;
        mem_ras_n       : out    vl_logic;
        mem_cas_n       : out    vl_logic;
        mem_we_n        : out    vl_logic;
        mem_reset_n     : out    vl_logic;
        mem_dq          : inout  vl_logic_vector(31 downto 0);
        mem_dqs         : inout  vl_logic_vector(3 downto 0);
        mem_dqs_n       : inout  vl_logic_vector(3 downto 0);
        mem_odt         : out    vl_logic;
        mem_dm          : out    vl_logic_vector(3 downto 0);
        oct_rzqin       : in     vl_logic;
        hps_io_emac1_inst_TX_CLK: out    vl_logic;
        hps_io_emac1_inst_TXD0: out    vl_logic;
        hps_io_emac1_inst_TXD1: out    vl_logic;
        hps_io_emac1_inst_TXD2: out    vl_logic;
        hps_io_emac1_inst_TXD3: out    vl_logic;
        hps_io_emac1_inst_RXD0: in     vl_logic;
        hps_io_emac1_inst_MDIO: inout  vl_logic;
        hps_io_emac1_inst_MDC: out    vl_logic;
        hps_io_emac1_inst_RX_CTL: in     vl_logic;
        hps_io_emac1_inst_TX_CTL: out    vl_logic;
        hps_io_emac1_inst_RX_CLK: in     vl_logic;
        hps_io_emac1_inst_RXD1: in     vl_logic;
        hps_io_emac1_inst_RXD2: in     vl_logic;
        hps_io_emac1_inst_RXD3: in     vl_logic;
        hps_io_qspi_inst_IO0: inout  vl_logic;
        hps_io_qspi_inst_IO1: inout  vl_logic;
        hps_io_qspi_inst_IO2: inout  vl_logic;
        hps_io_qspi_inst_IO3: inout  vl_logic;
        hps_io_qspi_inst_SS0: out    vl_logic;
        hps_io_qspi_inst_CLK: out    vl_logic;
        hps_io_sdio_inst_CMD: inout  vl_logic;
        hps_io_sdio_inst_D0: inout  vl_logic;
        hps_io_sdio_inst_D1: inout  vl_logic;
        hps_io_sdio_inst_CLK: out    vl_logic;
        hps_io_sdio_inst_D2: inout  vl_logic;
        hps_io_sdio_inst_D3: inout  vl_logic;
        hps_io_usb1_inst_D0: inout  vl_logic;
        hps_io_usb1_inst_D1: inout  vl_logic;
        hps_io_usb1_inst_D2: inout  vl_logic;
        hps_io_usb1_inst_D3: inout  vl_logic;
        hps_io_usb1_inst_D4: inout  vl_logic;
        hps_io_usb1_inst_D5: inout  vl_logic;
        hps_io_usb1_inst_D6: inout  vl_logic;
        hps_io_usb1_inst_D7: inout  vl_logic;
        hps_io_usb1_inst_CLK: in     vl_logic;
        hps_io_usb1_inst_STP: out    vl_logic;
        hps_io_usb1_inst_DIR: in     vl_logic;
        hps_io_usb1_inst_NXT: in     vl_logic;
        hps_io_spim0_inst_CLK: out    vl_logic;
        hps_io_spim0_inst_MOSI: out    vl_logic;
        hps_io_spim0_inst_MISO: in     vl_logic;
        hps_io_spim0_inst_SS0: out    vl_logic;
        hps_io_spim1_inst_CLK: out    vl_logic;
        hps_io_spim1_inst_MOSI: out    vl_logic;
        hps_io_spim1_inst_MISO: in     vl_logic;
        hps_io_spim1_inst_SS0: out    vl_logic;
        hps_io_uart0_inst_RX: in     vl_logic;
        hps_io_uart0_inst_TX: out    vl_logic;
        hps_io_i2c1_inst_SDA: inout  vl_logic;
        hps_io_i2c1_inst_SCL: inout  vl_logic
    );
end lab3_hps_0_hps_io;
