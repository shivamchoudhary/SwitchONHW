module test(
        input logic clk,
        input logic [31:0] fifo_out1,fifo_out2,fifo_out3, //output of the RAMS
        );
)
