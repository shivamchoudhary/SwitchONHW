library verilog;
use verilog.vl_types.all;
entity SoCKit_Top is
    port(
        altera_reserved_tms: in     vl_logic;
        altera_reserved_tck: in     vl_logic;
        altera_reserved_tdi: in     vl_logic;
        altera_reserved_tdo: out    vl_logic;
        AUD_ADCDAT      : in     vl_logic;
        AUD_ADCLRCK     : out    vl_logic;
        AUD_BCLK        : out    vl_logic;
        AUD_DACDAT      : out    vl_logic;
        AUD_DACLRCK     : out    vl_logic;
        AUD_I2C_SCLK    : out    vl_logic;
        AUD_I2C_SDAT    : out    vl_logic;
        AUD_MUTE        : out    vl_logic;
        AUD_XCK         : out    vl_logic;
        FAN_CTRL        : out    vl_logic;
        HSMC_CLKIN_n    : in     vl_logic_vector(2 downto 1);
        HSMC_CLKIN_p    : in     vl_logic_vector(2 downto 1);
        HSMC_CLKOUT_n   : out    vl_logic_vector(2 downto 1);
        HSMC_CLKOUT_p   : out    vl_logic_vector(2 downto 1);
        HSMC_CLK_IN0    : in     vl_logic;
        HSMC_CLK_OUT0   : out    vl_logic;
        HSMC_D          : out    vl_logic_vector(3 downto 0);
        HSMC_RX_n       : out    vl_logic_vector(16 downto 0);
        HSMC_RX_p       : out    vl_logic_vector(16 downto 0);
        HSMC_SCL        : out    vl_logic;
        HSMC_SDA        : out    vl_logic;
        HSMC_TX_n       : out    vl_logic_vector(16 downto 0);
        HSMC_TX_p       : out    vl_logic_vector(16 downto 0);
        IRDA_RXD        : in     vl_logic;
        KEY             : in     vl_logic_vector(3 downto 0);
        LED             : out    vl_logic_vector(3 downto 0);
        OSC_50_B3B      : in     vl_logic;
        OSC_50_B4A      : in     vl_logic;
        OSC_50_B5B      : in     vl_logic;
        OSC_50_B8A      : in     vl_logic;
        PCIE_PERST_n    : in     vl_logic;
        PCIE_WAKE_n     : in     vl_logic;
        RESET_n         : in     vl_logic;
        SI5338_SCL      : out    vl_logic;
        SI5338_SDA      : out    vl_logic;
        SW              : in     vl_logic_vector(3 downto 0);
        TEMP_CS_n       : out    vl_logic;
        TEMP_DIN        : out    vl_logic;
        TEMP_DOUT       : in     vl_logic;
        TEMP_SCLK       : out    vl_logic;
        USB_B2_CLK      : in     vl_logic;
        USB_B2_DATA     : out    vl_logic_vector(7 downto 0);
        USB_EMPTY       : out    vl_logic;
        USB_FULL        : out    vl_logic;
        USB_OE_n        : in     vl_logic;
        USB_RD_n        : in     vl_logic;
        USB_RESET_n     : in     vl_logic;
        USB_SCL         : out    vl_logic;
        USB_SDA         : out    vl_logic;
        USB_WR_n        : in     vl_logic;
        VGA_B           : out    vl_logic_vector(7 downto 0);
        VGA_BLANK_n     : out    vl_logic;
        VGA_CLK         : out    vl_logic;
        VGA_G           : out    vl_logic_vector(7 downto 0);
        VGA_HS          : out    vl_logic;
        VGA_R           : out    vl_logic_vector(7 downto 0);
        VGA_SYNC_n      : out    vl_logic;
        VGA_VS          : out    vl_logic;
        memory_mem_a    : out    vl_logic_vector(14 downto 0);
        memory_mem_ba   : out    vl_logic_vector(2 downto 0);
        memory_mem_ck   : out    vl_logic;
        memory_mem_ck_n : out    vl_logic;
        memory_mem_cke  : out    vl_logic;
        memory_mem_cs_n : out    vl_logic;
        memory_mem_ras_n: out    vl_logic;
        memory_mem_cas_n: out    vl_logic;
        memory_mem_we_n : out    vl_logic;
        memory_mem_reset_n: out    vl_logic;
        memory_mem_dq   : out    vl_logic_vector(31 downto 0);
        memory_mem_dqs  : out    vl_logic_vector(3 downto 0);
        memory_mem_dqs_n: out    vl_logic_vector(3 downto 0);
        memory_mem_odt  : out    vl_logic;
        memory_mem_dm   : out    vl_logic_vector(3 downto 0);
        memory_oct_rzqin: in     vl_logic;
        hps_io_hps_io_emac1_inst_TX_CLK: out    vl_logic;
        hps_io_hps_io_emac1_inst_TXD0: out    vl_logic;
        hps_io_hps_io_emac1_inst_TXD1: out    vl_logic;
        hps_io_hps_io_emac1_inst_TXD2: out    vl_logic;
        hps_io_hps_io_emac1_inst_TXD3: out    vl_logic;
        hps_io_hps_io_emac1_inst_RXD0: in     vl_logic;
        hps_io_hps_io_emac1_inst_MDIO: out    vl_logic;
        hps_io_hps_io_emac1_inst_MDC: out    vl_logic;
        hps_io_hps_io_emac1_inst_RX_CTL: in     vl_logic;
        hps_io_hps_io_emac1_inst_TX_CTL: out    vl_logic;
        hps_io_hps_io_emac1_inst_RX_CLK: in     vl_logic;
        hps_io_hps_io_emac1_inst_RXD1: in     vl_logic;
        hps_io_hps_io_emac1_inst_RXD2: in     vl_logic;
        hps_io_hps_io_emac1_inst_RXD3: in     vl_logic;
        hps_io_hps_io_qspi_inst_IO0: out    vl_logic;
        hps_io_hps_io_qspi_inst_IO1: out    vl_logic;
        hps_io_hps_io_qspi_inst_IO2: out    vl_logic;
        hps_io_hps_io_qspi_inst_IO3: out    vl_logic;
        hps_io_hps_io_qspi_inst_SS0: out    vl_logic;
        hps_io_hps_io_qspi_inst_CLK: out    vl_logic;
        hps_io_hps_io_sdio_inst_CMD: out    vl_logic;
        hps_io_hps_io_sdio_inst_D0: out    vl_logic;
        hps_io_hps_io_sdio_inst_D1: out    vl_logic;
        hps_io_hps_io_sdio_inst_CLK: out    vl_logic;
        hps_io_hps_io_sdio_inst_D2: out    vl_logic;
        hps_io_hps_io_sdio_inst_D3: out    vl_logic;
        hps_io_hps_io_usb1_inst_D0: out    vl_logic;
        hps_io_hps_io_usb1_inst_D1: out    vl_logic;
        hps_io_hps_io_usb1_inst_D2: out    vl_logic;
        hps_io_hps_io_usb1_inst_D3: out    vl_logic;
        hps_io_hps_io_usb1_inst_D4: out    vl_logic;
        hps_io_hps_io_usb1_inst_D5: out    vl_logic;
        hps_io_hps_io_usb1_inst_D6: out    vl_logic;
        hps_io_hps_io_usb1_inst_D7: out    vl_logic;
        hps_io_hps_io_usb1_inst_CLK: in     vl_logic;
        hps_io_hps_io_usb1_inst_STP: out    vl_logic;
        hps_io_hps_io_usb1_inst_DIR: in     vl_logic;
        hps_io_hps_io_usb1_inst_NXT: in     vl_logic;
        hps_io_hps_io_spim0_inst_CLK: out    vl_logic;
        hps_io_hps_io_spim0_inst_MOSI: out    vl_logic;
        hps_io_hps_io_spim0_inst_MISO: in     vl_logic;
        hps_io_hps_io_spim0_inst_SS0: out    vl_logic;
        hps_io_hps_io_spim1_inst_CLK: out    vl_logic;
        hps_io_hps_io_spim1_inst_MOSI: out    vl_logic;
        hps_io_hps_io_spim1_inst_MISO: in     vl_logic;
        hps_io_hps_io_spim1_inst_SS0: out    vl_logic;
        hps_io_hps_io_uart0_inst_RX: in     vl_logic;
        hps_io_hps_io_uart0_inst_TX: out    vl_logic;
        hps_io_hps_io_i2c1_inst_SDA: out    vl_logic;
        hps_io_hps_io_i2c1_inst_SCL: out    vl_logic;
        hps_io_hps_io_gpio_inst_GPIO00: out    vl_logic
    );
end SoCKit_Top;
